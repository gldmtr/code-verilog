module adder(
	input A,
	input B,
	input CI,
	output S,
	output CO
);
	parameter n = 8;
	
endmodule
